module axi_lite_interface #(
    parameter C_S_AXI_LITE_DATA_WIDTH = 32,
    parameter C_S_AXI_LITE_ADDR_WIDTH = 6
)(
    input  wire clk,
    input  wire rst_n,

    // AXI-Lite Slave Ports (Connected with ml_accelerator_top)
    input  wire [C_S_AXI_LITE_ADDR_WIDTH-1:0]    s_axi_lite_awaddr,
    input  wire                                 s_axi_lite_awvalid,
    output wire                                 s_axi_lite_awready,
    input  wire [C_S_AXI_LITE_DATA_WIDTH-1:0]    s_axi_lite_wdata,
    input  wire                                 s_axi_lite_wvalid,
    output wire                                 s_axi_lite_wready,
    output wire [1:0]                           s_axi_lite_bresp,
    output wire                                 s_axi_lite_bvalid,
    input  wire                                 s_axi_lite_bready,
    input  wire [C_S_AXI_LITE_ADDR_WIDTH-1:0]    s_axi_lite_araddr,
    input  wire                                 s_axi_lite_arvalid,
    output wire                                 s_axi_lite_arready,
    output wire [C_S_AXI_LITE_DATA_WIDTH-1:0]    s_axi_lite_rdata,
    output wire [1:0]                           s_axi_lite_rresp,
    output wire                                 s_axi_lite_rvalid,
    input  wire                                 s_axi_lite_rready,

    // Outputs to update internal registers in ml_accelerator_top
    output reg [C_S_AXI_LITE_DATA_WIDTH-1:0] control_reg_wdata,
    output reg [C_S_AXI_LITE_DATA_WIDTH-1:0] wgt_base_addr_reg_wdata,
    output reg [C_S_AXI_LITE_DATA_WIDTH-1:0] wgt_size_reg_wdata,
    output reg [C_S_AXI_LITE_DATA_WIDTH-1:0] input_base_addr_reg_wdata,
    output reg [C_S_AXI_LITE_DATA_WIDTH-1:0] input_size_reg_wdata,
    output reg [C_S_AXI_LITE_DATA_WIDTH-1:0] output_base_addr_reg_wdata,
    output reg [C_S_AXI_LITE_DATA_WIDTH-1:0] output_size_reg_wdata,
    output reg [C_S_AXI_LITE_DATA_WIDTH-1:0] op_code_reg_wdata,
    output reg [C_S_AXI_LITE_DATA_WIDTH-1:0] op_params_reg_0_wdata,
    output reg [C_S_AXI_LITE_DATA_WIDTH-1:0] op_params_reg_1_wdata,

    // Input from ml_accelerator_top for CPU to read
    input  wire [C_S_AXI_LITE_DATA_WIDTH-1:0] status_reg_rdata
);
    // ... Full AXI-Lite FSM and register write/read logic here ...
    // This part is boilerplate and would be extensive.
    // It would connect the s_axi_lite_wdata to the _wdata outputs
    // based on s_axi_lite_awaddr, and connect s_axi_lite_rdata
    // from the status_reg_rdata input based on s_axi_lite_araddr.

    // Dummy assignments for compilation
    assign s_axi_lite_awready = 1'b1;
    assign s_axi_lite_wready = 1'b1;
    assign s_axi_lite_bresp = 2'b00; // OKAY
    assign s_axi_lite_bvalid = s_axi_lite_wvalid;
    assign s_axi_lite_arready = 1'b1;
    assign s_axi_lite_rdata = status_reg_rdata; // Simplistic
    assign s_axi_lite_rresp = 2'b00; // OKAY
    assign s_axi_lite_rvalid = s_axi_lite_arvalid;

    always @(posedge clk) begin
        if (!rst_n) begin
            control_reg_wdata <= 32'b0;
            wgt_base_addr_reg_wdata <= 32'b0;
            wgt_size_reg_wdata <= 32'b0;
            input_base_addr_reg_wdata <= 32'b0;
            input_size_reg_wdata <= 32'b0;
            output_base_addr_reg_wdata <= 32'b0;
            output_size_reg_wdata <= 32'b0;
            op_code_reg_wdata <= 32'b0;
            op_params_reg_0_wdata <= 32'b0;
            op_params_reg_1_wdata <= 32'b0;
        end else if (s_axi_lite_awvalid && s_axi_lite_wvalid) begin
            case (s_axi_lite_awaddr)
                ADDR_CONTROL_REG:      control_reg_wdata     <= s_axi_lite_wdata;
                ADDR_WGT_BASE_ADDR:    wgt_base_addr_reg_wdata <= s_axi_lite_wdata;
                ADDR_WGT_SIZE:         wgt_size_reg_wdata    <= s_axi_lite_wdata;
                ADDR_INPUT_BASE_ADDR:  input_base_addr_reg_wdata <= s_axi_lite_wdata;
                ADDR_INPUT_SIZE:       input_size_reg_wdata  <= s_axi_lite_wdata;
                ADDR_OUTPUT_BASE_ADDR: output_base_addr_reg_wdata <= s_axi_lite_wdata;
                ADDR_OUTPUT_SIZE:      output_size_reg_wdata <= s_axi_lite_wdata;
                ADDR_OP_CODE_REG:      op_code_reg_wdata     <= s_axi_lite_wdata;
                ADDR_OP_PARAMS_REG_0:  op_params_reg_0_wdata <= s_axi_lite_wdata;
                ADDR_OP_PARAMS_REG_1:  op_params_reg_1_wdata <= s_axi_lite_wdata;
                default: ; // Do nothing for invalid address
            endcase
        end
    end
endmodule
